//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ap2Ms7wsLjlhAWg6sgr7Tz1rt873jgkRTWFFWWIj6i3WaH+Acx/UStT2Q7yQTQ3c
+lW6NwO313XugGilXNuOa8hAkgQGwRmWpE+B9Dw3CXO1ie9DfuKEFidRIVjsugFi
GoMbLFSMh3Ufc92QbXECwIlWXmUBa0gOG97SparTb/mwFyz8eqa4hw==
//pragma protect end_key_block
//pragma protect digest_block
KZms0U4c4fiH06G2BY1HuTH4mgE=
//pragma protect end_digest_block
//pragma protect data_block
lA9IbV3b2Bvp2iOIDs2Kua3fFnABdz/x7cRVJkC6oJNbwDyMP9k+AD6hWv/oGzJk
my0mEPY7r5byhXCXm4d+7qVHpHqAG3jNa/vUR21S8afXVOtG8QsRMai3Q6zLMsxI
VqBu+/Ne8teQtm7Myz5NyPncv2D2E/q+5qt+avtN+kADptgKnUOgKK24lvmZSW+2
hZA0pyA6PAsaIzud5wxBLcr/4nsRO6upob6r0okOrorBP9hb65MK8SSFVXChf1r+
7CCm2cFmdqbtc/yvxbJYmurTt8r/pL3IbV0tHe6WOuzXrnlV9dlvTknZtg5WQxiy
N0QIcR1PavoxsYei8FIR7dJ4ooBoQKHJd1KagIrmeu3ftaUmdpq26ZdTwkr07+v6
haPisr2n/JpgZ8Ot4Ck23zSEoCvI6ALhPoo4ngz5NT9B+VMNe52x6D2xZN/Qza2Q

//pragma protect end_data_block
//pragma protect digest_block
mNdvsW8n6G3c5mJSnrhQe5S166A=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bepIJpShuR3eBKETMzI7mgtWmkiG0GW4muaRs8XS8HggMYcpjZF8inTOPckR/VV5
+5t+yMlvDStqF7hLEgj4xRA7C3CbZKDqUq5WzFn7KF5XmBimacRZJfgsOYvIJhm+
E4lQQwYqg+OqchtfdIXrL80DbGI4kXTIKNuyX7F8hW4MgyypkrNt3w==
//pragma protect end_key_block
//pragma protect digest_block
eBTFiCZymfWUOoC36CwH2oACwZ0=
//pragma protect end_digest_block
//pragma protect data_block
/lZ/7tAAsIvACPenuCh4hT4OrmfePAfw5quy3FjZYB5JmKkMxVNvcwVSsQoudNM1
MTq6g5C9pR8Rv2n4gGyvg0bFyFwP7TuvoPAa+TiOsWd7FWKma2sDV/XSJd6zngJF
nDo5zwcz7i+Q6a9eVCmVntR4z8pvwxX0S0CPJGzG3LITAAVTbViXNgfE6MbXtCt6
U2M52mrfk2BoVo2ez6ZoEXpqDbPoCp2cOJ84Fee1/J88T8jP38bmt0mLZuWPE1XG
7IxXC6DsYDKNzX+eb+s4A3qVxPPD/8Y61K7GmrdPNuH1QUGDgli41q8V9tcQTuMO
F1UD/eE5flj9pVBqDXnTIA==
//pragma protect end_data_block
//pragma protect digest_block
PjqE9Kh4Uctdj4f5GKgZ0P9RAz0=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KJ8TGx9zGCt1ArVmyqpXTqjmDtl8ZNano2xo0rm4B5VVp0XRYoaa8BhiJ2LDs9lY
ezMs2szAeom2tY3FvOHyYPtwmPNbI0rKQBxO4DOIIfUPkrH0zPjf7FFB8QBLLMf6
EdDr/z7toKp/JxypvJ01FJoi77ZECPi4wRPry1TtxnCLFs4iBX2wNw==
//pragma protect end_key_block
//pragma protect digest_block
CH70P8LOw7vbLWWAGF8/SLig9ro=
//pragma protect end_digest_block
//pragma protect data_block
yboUzS3RL44hIdKX+QB489OuPgk1dcQMd0NIOyW95e9KD3pr/0zH/hvrk3U6ytP3
zHcHSwQCV8y3oTF6ZKsgflH9GibUEbETgEe/JpmD/MafzXwnajcPnBhybP7XyIyk
+AzQsDQgnktScFGTimhWZIZfMgnZXB+P3nNJCzoR2VJKFOfVlXQvlvP+AHuDqLop
RXc/bU6Hlo6W3pZkBhS2ccee7ZbMogTEHv95jJ7zWSiiwjoALnjpYJt1YoA3+WVZ
m3pv0XjbYOUBbg46WM5JhEK+zmm50v5NT5AUUpCl8CRQUR5d1Vc/t5glX5O3U1Ur
laA2rWZs5EdbM605lwL6rLrReWzQ2K2hNXshkXXnKA7XxK0/QdHazanNf4eNHnPs
QtxJju7fva0FvzAqUbhlfvg86y/tBb5zP+5tWmU4uF1Pb1RtYi1eJ5Kw7G0lA9r2
rnIJf6gZkNNiD23GT9fqH6ATY46ox98b/cRMPG8rT602qEEQQvYuNUg4XV+4003F
U6qJSLe7g1TJM0y/kPeM/OA42pXyvU7pVed7o1AcRvRQOM82EJVZB/k6AVjXC/fT
BxRTReenSj1Y9MDcRg3mAIRb3xGJMVlOo0BFluklViy8k1qYX4lyj0WfuRus6OB7
1rrDPdfpBSke7IhqpJH0Z+pKyb3sEsjW2TXHHel323jw8Wn2xy6ITeuOfKyJSaG2
3rQ+Rl+hB3hb6NYUi2JvoPrCmp3Yzup4S9i+44ZG59J3sOiRdKfKLyjbzEytfJcw
iHcAmwkQBNKcBdRQlVbMIKc3UwAcEjlRflHSRaJDTFObOQzGheh5DaHgWFYdFqGw
1++kr81v5lN7WA+Ljk5deAkZZPfUIsZsE2W6GTpdo1TL4+vdrUaXqRQWj4FP4RKR
IFgDRgEcOTAXFxWz7p8SluWkXFI+IIayLiEGFMbgJVQhAIFhhfITE47A627F9Ael
Onsv1F3+VOyqdnAhOsvbbifIl0y0IBD7VWLtyqBrlAQq0ddqmOine4Bu/xBpUiJy
0i98g6QDTfivVwdXLLkQsQkTLiYvqV/TWZj+z5E8RhrTljpdhHb0KyiJyVNvrEya
O3yFmW74dM8F6xl3vWclQcuPjnL0dxDzOBnNIIhdSuli1A52llyHV5xisMnPpU2L
Gc/UHEpLsVz8dygp7w/zcBIN/TkBddws4dWQJZpKh9jDUPfExphwUY7ol44NKo/J
QB5SJD0T5M39Uv3wzBKMV0T9TrxJskMaLxyyv6XA7jZ7Gu8/epVN+7fylCprwNZG
NNyWiIOoEDgQX39kOg88E3BwnPFaHP4s7gjnN5IsfPYwwrF9v+8CmuE3kbDcTKpP
o5tnlyRJB5XKswbEIHXMT04y/VbB81hBOHTQY/x2nYbDC8hatDQhb+wG0H1HLk7Y
27nqvCVMYcIF7wWQ4oD9A71GUcEyzZm5F7m+vKg0rExw49j88IYPN3Wmq2xK+GgP
HzQC942eF0M3x3pIlUafjIbS4NVZYOd4W3jL+k1vQOCq0C8fs0s4Ah5QIFXMlv+A
1OSCZ71DlhNLyi+iStI3VzEtVJXXMeu3dtTZbq3+QL/j45B5wfUPynT2Cy7MAj7+
zZnYc1OHSHx0MB6OvbwRF/sTW/Cop94DhjE5oxWd+8MyAIWTw63czkJBsWzkRvE4
cTwaO9rRt3Sy9EojOnMtd7dxni+kkHTNbLY+jugRfsxgU4lnOAlXgcuj3SxmacV/
efOLXYI9O4K08b04xZZCYeVgY7iwxNsQlXGzni3sQjnnH1q/6FQe0qrLypHuxqK4
+AGYf1Sszf+dJaxJbIGINAi4ezCOtYuMEuZ5/0JDzNqxPcO2TxW9MmSVtnhMmDvH
454GCUIlcmmcNjDCbhnIG7xWHgiP1r+ASbjVY9rz9Y8sP43UUcdaQhBPlUI/P0i2
rpoOaJllCiF/csDwsxyl339UwPOLG+yGyu9gONVa4q0U3b5GpM0K01Sv7J0gQI1F
1FKUF8kqSY+8xeVpxROPI+HAt6lxt98I1DI9eZ3YCiOBgdeFuxjtqDQUSr9hD4n5
bNWW3rbSqWDKkzknHXmb8sNMRM5iSONeQ3BXeD01nd50cfuA0llwRz7ptcAInnDI
w8g+sWI7u7gR9MdzzCk7Y1s2TGpz1nmLcQhs7qZB4A5W8DfrX0PeoNp4g9v5X/MH
5TYZS+pC+NaECT8Ir4U/UTj6W6j1ktdDn1DroCGr16EhW2XK7jpjCPX7Ln2iPJDM
p1qsPHbv6cqKW39tvTNBNBga2SrjO3CPvRcUrF55ta9+peEmFwzs7aUmtnSOLX7K
SY/ckSl5KqA3mdXGb0uUZC9Y1qMsI8eFtskVur1KR0ClJYvBujM2RiOg+vPDiaOK
QDUJxK6lO8ssI6zSUfKLHJ6QaXv57FlzKDzHPbYOecCRKCnjANENV3sn+y2Y5V68
+aQoSx1OUyidJMXBYvC8y0uJsNfsjWRsWeuHFnZ/czTds76UE3C5B8olPYSdDNLg
Ce2lKuzDcB5YiUAhusJDBILRS2KoGAR2mIrK5AtBRVzAmrtwFTMbm46StiIRXB4q
z4OPHsoKjxzmWr7+r4xVmAsi9HLJBJNtGRYdT0hydokWeBbk6vQOXUUWi4c7UhVz
eCnW4zMzt91x9U4/bsVuhORFPXzCDbjL/nfSsToTr4Zx3I61ilBW89kC2NgwRzq4
dAl7cuNRyfMVYz8JShtV5vk5PuT7GpZaHTAAnch+q9XXsT2wW0r31oKHdW+MQm36
/D1mAC8zgKOvopQb39O+F9iS0xMZmJQNNnQFKEjNpVy2WTjedZTsIe4LT7XW375h
N2ZWdGu80jrI9Kqsne5vlr/zoLFuRmMYjMJOUVFFtyQ2/mqSC0M0W1PhdheDziB2
FVxM5UugveY5LOk1R+twijMkd7llVdNnmdxOCPY4WrEuo3FFm6f3W/mUFU97x+GS
LBgRGZdCRNGC+uYxng5Kqpjdk2lIjayU/Yxv4vNYX+0vrprm+XduBJzp5zBW0DpK
5n8KkNNZA+mph641N6KkRg8F+j+PzYT2+km5+oNA1cDrrJe6VWcoDyLo4G6Ku4cm
H0s7frAidj29u0TMLxQ/7UcZGIuE3ALK2pl9xN7qEgS2uH79q1gv1DGTjWs2PRFU
9KZbGTDxm33X/OFSDJz+0+fhTGBwVaxQFFNRr6gwyNLVD2HMI1lksjZ/aawhElN0
xFPj7iAQmcrZNF/7G+awjwPR4sRZPTNyA4QZPewRisUO954c7iZW5Fd1Hda/otOE
g/OwrAIBLrvUHsAIBrLM1xzdPdnVigJZhf5zR5/yjCiDpsd0GyTQDY/LFNQVhHF/
pYvoibEfSbdMUnIProTar+rOiP3ZfeTCqED30mwVJvODWO1SRU6Q99MVxMEaODCs
sY6bbp01C4NIiTfxnduDbjQp1o+BlywLsFOkchTsZn5IZmgMVfGNQqzjuuu61c3P
pq5gdIAXpnV2zKeyxCvmJxCrH97KN2muhYhWzzfLDVT1dEYEhuPLCtJFop2OA7cO
KgYtCkHb8WbuIt/rDnD/Y2+1djtM6/2qYyK6QbxLSitmfnlzWWByyd5qEZQJLkHA
IAxHx2EPvZUsdSrFXam5vqtTsJirV8TUExPx/C7O3kaZbH/M4PlLvGNyqUa32jTL
3vy++jAAjeAY30d6KAfI2if9QioqFdb9tezJIpvGzZSNDVNVpVYLK/c41jpL8nQk
9o4OrbHdz/BgNxSC4WGl4FF+16cxE/S5GzBmttfDmdxu+ozs/grTHh4vTIGryBmA
+LhGJ0oT8Y1058UVJtLjTmoZqi+PIEwZPYH0odtZYaFl3MKfs2otMubFxXHZMJke
6b0Inj607sI8OaMyIBTw71cbcHd/bh5pDp1XW6Y0TvkYmPh+3DjBQsxtw5AvahMq
74TMzWbOmck4lkk7pLiGdyzdsisk58TSc1kQVXrKRpleNf+mZXKQrKvm9Ta3WN4S
01idc4hVvQ5MUEy0WtWYm54Q9bpuA9WJuxAUq/sTEDdg+G6LuXdpTGxSvxVk8M6L
2MUuKUteyxdzrDSLgt7CsNzWni9B0YQo7WJZt65nCJ0n4xTNSdOYcI/Tqdxjcd5O
fMB0FhfM4sv2Sp+CJ9eXeRH9Tw4YS3wSc7ZPuaZZcdOw/JQjuuGwuoeTC/tzEbgV
gR+Nji530cIrnnLqVIUjYtRjzcqeBeBgrJ4Y3EG+lIcKr1kAkOxv0VLLUuMaEKQf
eg4x73neIVFtp6nge54H08pE7Qf0DZwM6f2EJC0YHChRLunAYRfbvu8DC+19Fw8h
Mj7nE1DaXMvR86MoI+fbstodJ6st1MIEhvZg0PGTA9cqDy5Izzwg9HFGz0FsD3T+
UwqfHpFGWnry8G3YNwElVWjHWex7QMe538OuRwcAGTw7jeZdf0MZuTNiSE98oCxv
TNJliSm8Ruz13dVFyroK6rcidoPZpjT8vASCQXj707ITkoaMQCG/bB/D8rfskClh
MLR4JZ4OpnPeyHXu9bkWu1Hj86D5ecxHX3JisoM18n6P3fSFB2Ao3tYdRawmzA5w
0VwGoD380YZBajXNpvgMZn7Ko+MEqsex2NkF+f8BY9Pv0yQqDhkv6UoORQADOd/M
lZNhZrUnO6IEI1SNNo7/V10mt0kWiaQLURNWpfQw8h9LJCiD4NH0N/axSFtYGXJC
tmUAhqBF/7QnlfRL6QW4XUTrEeE9gfmYp8CnDowRUWWUEtOIsiofDeTT1vaYmGks
JFRSOnklVcqw+2OEjXNV7A7TMrf21DXrN7Fkw91r+7xy8A3+CzBC6LRziQSPWZNS
mn4PYXQUURhA0B+wvDBs3nzf8RW+jfziDRrZ8a0ltLKiZnHwwAktdxJocGitINZv
lLWizEcMUDqzldpJ8M38G0ZA7YZlmndb3vkRQn9/2VdWGLtXOiEywB9M4uLVCv3W
3SIP4IsH/96InGHTpooh3MXUIZ8kbJEQZoBTm/FTZjedG14uqrMDxsOaoPpwIe7N
9rNP0WTvM2ErsTIYfz8I/LT3mttfkpNrjZUXJbP7mmqML73jxayPRbMY5cTOMuis
3azHzAVyqkLRppiPBmJmrciNwiFjzFYKDJrTJ39AbD9Eb+DJC6hXhSFMARBChUaF
fuMMai97GHikNiOefLCfH/EsrCg9fo++Y0gNiRYqBh4eddx7eUWvDUtiPlyDCwfV
sN0Hyl6s+jB2Fh5rzo/pRtiDbeTrMuMMKHGXYUu+S9PjtsigUNBi0yl5LnbvQ/ny
McWgp9gbp4hFYikegsoSRTi5oBM0j4fofw7Gr3XqQRYOeosPwsiS6FvBCOheEn8Z
MonB1YGqpTOjV5GCe03kSa4gHZgER/QCwgPLcnMcYbuR/qY2sCxKzkIt47BUgi0b
yJ5W4unAEebjOAxYpaTCtL4bXfm9Dw0ta5DSGkXw1caFLLV/9ejH8Xlv+vJTXPK9
1g6lC4HyBspCO/pFiiZTLCn1hchNhTBi+9EFsWO21CleRV1HFz3GS9W3QWPnvJYC
T6Fvy0YZ5K1BuThwXVcvAngri4FYh4O//DbKBdMkOB29YWPTY6x9C6MG58hAdqDv
3TaasQ0R1Yqvj4HqBIDAHYqh8uvImQupDjYklrBO8NYPQv/m9/fLKCZz0mp4bULg
HudGbMsACwq9w0OStlCrhufrCCRoyutUn/4miFvi58WFaui014Wvme4LP/Exw7tt
29y0SoL/E/fKcw+Va+NnSlictsQ+XLS7mr5XsqWDiVp0OLZay8JQ0hxA7sQBuXhk
zqHsHdrznwNsGkg4IYu4qb9C+JRoIWq3oDy71vhdPQpMpHC4n53/9ZGtNow+CwDa
LZ11mcv8/IRzrzhWTik7xI8If14X8yLwSmUqtGON74Vx1Gl9slygEKKRf9eWbWo2
yUwES1qcDWBlU2ZUf0uJFz7L6gs4cuCtZAE3eSOvDtM1nj2bLZ7X96irHW8I9upe
4cLAyZEffItqjHf6RjzV9IS3dmj91Y0tETW7sG9mWf7hU0jTFK84Rl5gb6wYDdnU
iKNWuFVgjSaBKu0wC8sZQNLQPuSpX0h5wlQiM0N+carvYiHbL3l0fCvogoKbatU3
4f0FO0Fu+CnsOmrsVZKez23FMzWAh2v6BxytVORfqw4k6YOj1igdXMy/lNKpnSI/
f5kQChq0mKW3f/1AY7sPAgUk0H0f+Q3TlXdOTVutulzXSIdN5q0Vug9xX+Afc0Ek
jsM4XQ+O8z942v3OluTdy/+eUNg8AnSM1GMS+5gkxOD9D242tg2dlYGbqZ+fEYBo
EUcS69qf3V0YJsByP4bHrP3ge3WWGTDhwxeznEPmY7Sq2TFeaq631ZPubk9smhVc
F6MWiW8sALpg90Fb743xww6R6m9BEdiAUC33Mr2tWvpRSJICfk+VpqrTC8aZ8dbX
q9hUUrPnIQugQMiGF2YU9v2Cfk8NZvpmLHkJ4Q6kmKN1xuNZtVIehqhkFMQK4R8D
MGpiBzVhC3TtRU9opNnSD0nC3jE4lGisj1vmwESfhFPYipK7ykMiWH+f2OM5vbCN
X0LOKeooLdvRAd6ZXMgAK21w812Sya4GTp9f/W4iXIe81raa2tQA6Lgcw/h0jM09
fT+C4PnVKgy9j5M2NKF0thGBMqKwYOL6CYc6x9l6ICsO2grUcaB1XGvAV+/CDnzr
+zGU04ReoWScaOpd/GXssFKRV2YS12HePck8wYwc55tBAh5AYp3aZm/0dPehTt8A
FGotU1U1gZ22Nx53Ix+/g23ej+u7vChnl0h1hRtE3YZ+dDezh/8nrBMQbacYnsCu
OkG9ESdHEnMYnNrnaRYRVzS0keBoLR7gkaXdOD231ZT6iEeR4fmymhi3j27Tvd4R
TxLgMYKzC8jkKZccI4L54d/c8HBq0iTa7KanjdKBsu88Y9Gy8XYxwGt9DxoQbuzV
T3Tzm0xpsb2l5L85nDfwoLm/5lKwcoF3eDXZKLA28+MKUaOQH4ClI4//OX1KUGnC
YoAbBsH5y6TBiHtyEMS2G7iRjQHcLA/Fdlo0nIi9gZb0ePiKXEUs9GW7G/pN6TxP
F3JddgEpx8FdRbpZkI6bEawhwCMgkcSce+I1SwsSGh5gXeBhXYX7n6Q0QuydIjbU
uvE3SO2XW9sciPeEI0PozPY2av2uBnUpt4qoSuLdkDefSh+DZiwrXC1JqFTKdTVF
LDOEBR6Dzf5xHVnlMOgnhtiBPWXDlnAbeh7OwJn1RX1RGgAij+ZSrcDZSgFAZ7DB
kuFFXLoI+hzAvGOpnj1jj0lJ4NBHCaryPBx2yPfujr43MkbklDCdgxMZVfILCEe4
x7KrNJtvimflfcya6mW9OJcVz4YgGhFwbdl8E+5EvSQYsutmne0U9V2wNKEW7hu0
oG4Tyo44Ua73M/5z/s6fFZKPJ6yyI3bkWI8TlFViM9UHURyABEAtVVOFkuLYN5VK
2msEMyW1v0AVqbEbtQHMvPgM2jjEE0RU6nmTB+Ajdk51o+d1dR7oUQQSlP3G7+kX
OCFqVDFROdj2r0g6F8tA3CE4skk6IIY6yKudF8wx9p9WC+qODpV990Oznt6v12k0
TtvKgtVmIFzFsjBCQmZA4roWOtJMs8aLqwAqOL4kzHZn/dP7hmSFQrYMPGP1XsIT
EEKA8WSrSHzQ+4SjQ6+rHuJJ5XW/mVXsf9ebL+rtKBFWSBBMqPVccKk8jItZh0Q6
8fdBpY1oDw9rJEUZ3n64DFnVmKuER6K/N2h3qNxFlzDUAgBm+CKuqU12xa+2f9ju
XF3oj+tuRRArvpS9v/X3r+5ty3gIbAy1u5ItaCCio0WDjNjXACbpMM8/uOOwNQuB
4bV4tsMqfjzlBwfBYEuBdY3RxvDNo+XRB19fGHwX70thWhfx9V8pjjBmxEd6E7ov
XqnnqsvLE2QSYqfiMCIURRh7QXB8Y5Cr4v8ljFIXbOOR3SxR3oU/hFqeWfxBJrrV
F+qEuZLasNc3W5hw831ge1m/l6EOJtasgUnfw0BbEW2L75S3Y2KK4w9wuxQnlzZp
syS0e2s3SJog9zfbZGVKysDJ+CEmERQIH3aFHAcpz+sJDhOXQ+i18bWwjMmUHTXB
4jG3rHKdDC52T/V9DXrJVdEODEd9MKDxcbEBNDU2DAChGs2VqZ4U9wfDg6twVYgA
HKEcc1zmT2tv3BTXTT/ImsV8DYs9OrMJQarVa1440JljlyNqg43wkHo4auhg3UsI
c1KJ+JANiKEDInaWD/v1U5BmkMgcc+pDXG3+r8csN09Y8rTX49ofYNVaLss5mDmm
BIBeSmfdhgy9gEoETQUdPhHCmJZFK1gjuSVNs2CWv8hhO2LwxMY2lIhREj4wPsq9
MvqBx2usDeHkFZy6T6fGq3PwvYt3OYuuOKDjfjd3n5uLyxEr79CJeAQYYHhFL+v0
yXXnSQ4aACx2+AAcnZLHLS7mahwFWjH7Ia34UFowyXQhX76NNRvqnSdgoaJ+Cc9D
7cqeLvVQl4pdTKKZSLd+26nrX0BS1G1NTuhAfx+jVcEnrKiMSfqmNH0RoeIsrp2F
srdcixCaJmPwOhWHWmk5F/3TjVzw5L6Ia2HxC2NDElA4EeQARd0vB2coeIylaa0T
3tsAeghRBfAPNBTo3s84kulmyDRJyMwdtKKZRChszA6NLpD8qo0naHAUy6JO/gCq
PNKkWOe/3QqJqVQZL38rsmbfxo4ePI6HmVGKPmhp9Y6dKUJzvStoYqUMhCl5hpiF
lOSUoDWiWdehsUqJNiIky89wdj+jmZ2nFesBsWEmIY3wK5oedeM2lMnzB618ZjKw
zrgA5CnWhFFL7cwMN9L/IDdZCKdgzIYwyOciaw5Z+NYhKGRS6ozQZjkWlD5QceGf
HwIkVnLWLZDPTliu85kQmxsukSRz3SJip/K/prmfYzsAvb/V11KgbvL45sCZYvb/
xuSeYu/olC6qmptfi2QZLDkiFq9nZtl6beRgACMXScvSl3G/PXpkHnv9vNmqELp+
pwx64oFcUXuqkwi5hF5fJ+q0WT1hnRT3So0oPFeZHEiNf5UPkNBpaa7Yx5J5ML9e
HSnvkMX2JCOtFNQtDzi3Wb9SA/9xsnFs54XNFFGFxHg3EE7OGSz1U2B+fIYt48ig
BdU/ZtuHf9BhYZ26RZHepbwRkZgjVmfcM2jl41+B0Icp31Y3IJEilvUhdZ+bLS8b
HHDmZpjRLE+kPqSDLHPGtArpgcIwqi63XRky/kDi3DR0IPQavi9AKQSnLcZOwCuX
f0pseLB5lk4U8qMOMttvuDBUGglEVBK1qkeOo014OJxqbYxn43XctPG4sRyMtV4z
wg6g3u5+DT4Gy6wXdDmtBYvLe6MxJE1bBtY4gZtPg/9GWtyelgWK3zDGpzK6EC5x
JfA8L4hKKZd8eUXv1e1o0M7USJI8XAHjx4Yn8RMjIVS6rtl+S//5tv077VTJfvYE
R4ffErKFgFrRoUWCuvjEHce4JHS+E2uw9XBPL4hwUS2tQJZUEv8LsY9thhN3YWzk
wtRoMOUzQHDprpcI/qc2/UPqwakIfiV9c3tQ4CNPOeanRIvISRAFIXl7CW1tzLLv
NtdlZY8+TdO4zW/GWppRLCD4I086uXnyLbEDkuhZwracHqAK9KRqut/kPKvTISgX
+tCisxoCUu5vnaVJ4A+v05RbBxTDgD9G3xR7LtHGjulIDI1S45+PMvWo9ir8yLYi
iWeaA14LpYyQcE5Z9wF/NFi0I6Ekj4uOv45L+Acwl43BaPuUNZSB5Du4Lvmkg5a0
oP1xGyqVjFyXWKjAa+B7JiHt/GpC0Nn2yav8eRFPVlQdLipA9Pa3F2s6R+KZQcOP
DyLSGCRsLGQBr17tqMkTNbKD4rozyA3CF2cgGAtrtxLbHi5xxAv4NB65CYwYxUJq
0fHaeDHfj48qOmaFAz+Yv5kgZJ8RkRxpFuI+qXtd4F4ZZPY5tXwrqKlodiIFChnG
9VrDZlThM1PPGUFKaqLQDkVhrpgB9x41ZL3nSvnfFgB/fovu+7K1zUeOn6gcwFQW
LohrXvOlGK+qRuiIYxsgWSdbPA5b2fuOtRsr48LUHVjhvEdBaWtZFbw5xZCkHK0u
PwEtshHRucZttdfrK1icNbvL/LOuaRYe/Tc4LitrVHEJzgQh7Jw1GEwd6pKAdgzP
eMjfLdahK5XHnklBoPq61+72lmznf0qY3nx8mc+fgVNRUnFTnEg+Lssm3GH7Hchy
S+BH42rSDeqb59Tc6TKOCedpUmExUfA1UnWNHCh+KquUQKM5Obm7MUrouFd/R/nE
QVQsB9QGGCVf23WwEquO5MnN4VweqUKGl8hc6jtQrCQl2p9MpVeO9Fb1C9qyYRE8
nHTTCpsR0vJ+iogYBQ2OLWj+Jgf9rLH8AxtGludrdwD5I9+gA/64BjdnHHK/jjFg
2dDWKDb5oL4zsqM11rXmTCKglKjgGkbGYwsoBt76X9KNf0RLKQSUNpg4cmkytU0G
7G2es9US/hBAHwDMmxEG0uV+uRMZhf6DVgXM3Q1Vb8lb6Xu5qs56yruUaSMx1QDq
gSuDVPu/TJHH5B2ae+e9quLPIhn/Ipg5908Lb1LT+LwtBFIb/ug34z5dEfldJ3bE
wVTiHn0pyuTGXvxfJKsP5GKBTeaj6y86mUz4xyRpE85/AskmuowTU/MCzJbMXlIG
lytkkxwt4f1ibbWLgU9/C6GsYqSvm2xI1s+RzTz1Gx0IohMssb7g1pbyyez0jT1V
dI0rCixahBpMXN8gtNXJnrxPrWgdYlzXJMR0oUG2KbeUyMWxgoLA1WVfaca9w6zi
weZ/MyF9CkvEVc/4ILCaqakVL/balpLbLe4qpRqut2qC4ebu9hxrjCM53UQOAZQD
KQRQtoOdrPK6/eI3SX2TReBxuYyx29sijCTXWH2HiSefWoHeZm+ASvlEBO5Y5+eV
3uvxjCggMjuMBs0577dmYUAMGnxKGU6PeingwLJw4OobXmWDdNJDTddULThtVa/4
oRL7tb6DQGIINeyDTrxsRdFoCDNobtddufGQJhpj/kD4LWQr2NQCDicmHBS652/r
oQWI4AKCmgoe73Fm1+9wfjjcFozIrHqKWtgjVrUEZKByXu/OVZtH9UiuJHDJKESS
RYwvN/jc54vjM2GJSTiRpievEXJ0eTmwKCBAXSZV/4ZDG0Sc+TMcmLka7wny+kJz
qKdbLj+/U7IqPpMixuDUDSeMKVwQT5vTTwYRGaAwZ+pb6IvzdtfMMC4+s/RNnr3d
vMxA1Qwao3L4fHds+wleCtLyyCwq4w3byzrG7Xf72NAt59KZiMCjEddb86UBTd8y
y19PqjwFZzPImjE9YMG8dAZaS5nlKfTgpoYAOB/Ff6liFyBmyiFZfPRmfRd5zy+I
q006Bmxgvb5u9LankB4zeeXhUf8bcFe6Aoq4qS0PhTSp+ro9IBihw+Qic6bXumP3
enNXJRwkEN9qSi7chMhAnWyYxS0tUkYaeieYPDv6ppQFU9Qy4fRKmbZH62nMdhMq
uzSr8mthvSjyeBGZG87k3hWXXET5feTYFItnk2vsZ8uDrE3d+sHb8/hudQCOHs/8
FC0WF+FKU3u+/pRyvpGqVCH0H9vG96Za+p5qKX8k2Yre/l6lYcDQk6JoLEaIG52i
SNVanQXRdIXvFQRjIDfQIbTNaT+gitz88TjEWNIOdDZ5czIBOUYYM9NVpp2MP7uf
2DNVkztIN9prUNDK6FAFPzJMHp49gbm4if9dNe5rqKY1siVGhgbAzAEMNjL06F+Y
AgnBuuTwDkJe7Ca6xaW3YFxheMskZZEK6JUCMRmHpn+82d4tkW1u1Fx7ld25TKJ1
7OEiluF7DWP0NNVqnn4bASMetYFwCs0LIvISWrcWUxgNrn4WleOtybWFWZQd7xrl
cmhlt1Y577a3Otqson9O/NE+NWzKcCvrL1L423v0I5W6Z0YM940r/lhRquJ34SGW
dmiZqk3njQDYKEd/jdZmpDYVUT4cp2eQl6OfhrDOXP9Kqmn3rQYwzIA97lV+HQIC
rzoPnUQTU4WK5tNqfUqGAxLkJMk8fsi/Ysf1Ce/fO/d5QwQ5jPabo82T+X4bthZw
VoCyEwcD0GOcShhSEJ97fOpQEdYte3HxjzodNHNHiFO8+e+G0SHGd5Iet2WP5uqg
r5zXd/BZ2JoTv0xYdNMPk2mXu6CV9udwyfdK/86N/9C5EZ+/B2D1wkvwpOhh41Fu
nfziWC5py6S90twbygs4w9lle+A40KgKcLYU74QCwT6R2ao29ATF8eCh5SUH+GV1
KUNJC9JIE2tAfwsumA58QQBKrxVuanhSHmufkBDUwFxMUiWMRz8R/+wBi/d/YlgB
W6cOPzml+nj3yP3yz0OSWwT9gaJIIzDO7q1DAKwmdsgnm9uoTrTwJAPDy/PYCDW1
D01Um0VHsVC24i/Mmap2tLFS1KYRDgtsE04x8X4zTiHlPEBKc60Y3PEW9KDfVykF
2v4LB+Pgch+TP22dZOuEBZVG1TCf+ZWT9KoLJ08NFV15iHPbLKPFxCYky3f5yKV+
8IT0DRIo4WgoFLFiVn9KNwlk2/ZwjnCAxgSX/yMMiiPZhlLFQTS7oDuRHIe492oU
2hd0EucWM+XTlEz5uj2Y4ae/vabDvQgavHfEIRApHPHnCj6FTUxth/MwP318VEvq
DN8vJ6tV2HPg0HE5Rast74ktGAugQ4xH7VztJeTDxoGcPEosbx2HAb+YPn7xL8vX
AnX8dIradBs5EZgQ0kUueDfccDNQV7y/u2GeE7I/loNysxNxvDi3sw0sw9boZ2X7
bu8hgI/u8Ni5NzcL4q23EUmKW0nZL6zVFnV9zbwaDwg/1quQl4j3AisC4tLJZWOC
jKbYsipc2qRJCE3Y9i39ee+5Xhj8SU4AEE0T+5NQ3cmHr5kSGP4PYClgidUnkXyt
SC89YgSdbKSwyzyb99mJttg0QsPwdfYP47cMqvQ4mfqNtcJpNWNkiWGRq6kOdk2B
Wx7zb6+HnypEZJxTmMKj1hr1SoMz3b21I+QkQV1m/Ruxcu48wQE/UtXb1JQzuio6
odP53K+3M1m9JfJiMS8wmuMcIsCCUEPvw1AzqoungwhRAB7kVijhM9Z1mxrw2/5B
djdvUM4goPd3pde5fIEkaFQs0y7WhtE+3dlQRhNZz93fDM9i0tMtmnIRBkpX+DAu
2FrdTKFQKS3A3TudDmb+vyWACiMh9YpTxYCuKqFjomqIBFCRiBlR1pKI+QqnOXSB
kHRz6zR4ehQzIvJ8YrdMJmqdZd5DvQmrjXlUqL0sVAz/b1Bjw5JoXEqWxyLtHSB4
yK/lZ8olmpCwYj2uJnL8bYSklKLcenhiuOPi+xVn96Ub6hISJ0swbIHJW5TeqG2G
OSc3ELmCO9P6EH9tH+dZ6DMX4AJy2bWrKIUh/fCZUQx05Bf2QQYBS7MLXXTOyDrS
niEhWddoLi6uAkiAkNANaNl/+j2/W6YUEunQUDLE0gvblznFiYA0DvO2o4qaVzaI
yzIvYbCtpf7JafXbb/OUnUk6Qdi4vR9nGV7KeujBN4/Hp9I7AxWzU2VxZZELoVPR
5hoPnOtwK2Z+W9Q2Z9F/QQ7o4UaUWcRBCTA0SsnMtzSVCYq5+XJ9yUA2l69u6oiP
c00BxwGsYdUkLmh0/EV03D7Knt+soCKZUzlhirC5woGAqNfAUGMX/jNKzBghLIxH
/Em5ue5rqpQILBqHHRzMYl2IvHPA24A3ZWKQ1eNMTTY1ZqyLs2BVoIVy6+kBauwo
J4XCEeCQrMi5z5WnP3LiPgJkiqfK9Um+p0hb7ymtxvMy434XkqSepkL5qpTgYYvY
SqpN0AJ1p7mrVW9BeZHXh8lyBjMbiDUBjVFuVNe/RtiBQ12A2PGODXdMgo5RO/Rs
7OP1nolHV6dZfLpKfbAdTE5Txe1Lo6uxQpJDv/rXEa3sZ9cZeNUN6YM9avBT6krM
UgUfjV89Gn+7Y3GarRsgtbBagfS4fWKW0Q/Frao8PaHokRuH+W5cQu4NWEp63613
0gHpe4Yrjoj+Pco7Wza4K7LaYa6ddtoNmviAzJyuiMDrXLI46hdNJZYxIrhQ5uFx
oHCnDNC231N9Y1MS9cs/Eh//NstQimDQeqCM995o56laXzxa6MzuK5dl4c6hl2Ji
d9/ErGGCuJvbX5EMVdfgV9QZZzZLVHiETWVISbYBdDfJQNregCda0O0UJYxbgNTb
zl+pO3myH3+FlvuTFQ1vRBDUk6U/i76YI3NebBJE3zYouMV3hzmq0D0X4QYS75pr
Mr0mU/eu2xTThgUgANgQrs/E9m6GO3eyJa7r6C/xWkTHYB7/flRjZeGBlnJ8tVCw
clNuYhsTTeYefhzW8UpGsBNbRZXnzyOo6vtYx2bunyUte3JwNnYP6qnUBgA7tpO7
wnNsmBGuoGtMV8qCay9RSFGesJ/8DdVC8Rs2hH2mGXDvEqYrqSfvyvwf8VR7AJBm
4yjwqffKsflratm6KgzFuRfGguOfAYgIKSQIa+OaEyi2bAw+nBIiTYHxsMq7s2Ew
E4JaMS1mzpPvxUonoLeCTzpxnUALigFF9e45J4+jKjK+lCxY0A2yHm5IkQCBN4/d
Z/+8szTuaJYxdBghUPEymUPPUlIsfeY9s3vs6rJY6J6e8+5VhZ3zLbug+vLiIoSN
FeJLe6zdZjOdxhwElH5vjV2shpCK3LZufPx+AULr527Gw4Th+ml4QYw0Sy8rf69j
lbLP62oBOa/u4iW8uYv4002Jxwm6L9n5bbwAM4E3gN6D933BFzJoeW3rqto0yNYB
WkvlKftX27WJY26h5RZL6OcafdgRJ0FzErtFTez4sVsFp7EwC0HA2FL2Wk200L7y
MfZBG/V78SvVPQiw7j9r8/IPHF5F+XLhtOFHW5MUSrJtwRbQW5nIbEuc/964esGA
ChLQQ9XId6Geg8T1CC13TqmI9FbooR3GTra55mSr5y+ekJYq3v8Xg/GVyGeTWIFD
JpC/ThUC/K/y2NF4zvUmtlD+ndhYb1pyzKpirgONMtxTjMmqIYY+0vqBS8jSzBwU
gXupNMOAEZXsu6NsEmLqVJyTjHifJZhONyCM45bNp6p77pvcbFPamqVJ1ScXpAMp
DlccATMlbQxkERznayIDybySPSX9EVvJWu/CIC7dYzCOgYnkIY77Zgt9mK8GYnwG
nGOtLrFe154Fond+gG5jMd1LIvIOuFsipLARnd7cljXINRalgOQ2lTxQridj6TxY
TIMSqwMrXUyB7gZtIoXl/mer9RoeF5BB08iaAIw9PCEmqO6hywnMGQ/JJkIhgwDb
sTY3jOL1R2zm4WIWmKoeRroX3chiuwDUrAlflYw3r/Xg1i46AMMbFGCqaqfieRy7
e9TgC0b8tlm6gU9QvReYRf9n13N/newc+IGQGuIBrO34bPKzDOBoBTIOQc1N2dCM
F31PN/JWJHLkZN4a79j2v1YtM6DMhzs6W7abR18rk1zamjz1NiKUO+StCdbEWulx
boCAwyIJwu9qGGXr8XEDRJ71eYLo2fA6yGNJGNY/albgM0OwiBUNHHkO+d9lTsho
J+Z4KY+IVVvWn2goFMIFJb9AA6QXillrASnH3qArg+rLKabLAj9SxBLARgTCN64L
yabmbu4T8tllmieLnZ/IpzQPcrhnHF8X9PWo/PpNNdvDl4bSTQSACaRQAHAGiItN
aJM15LeGQMJ205x1AQqP8Z4wOShxsYwTArzFzrDguQBNI+eRe9xsf7inmdHKLQL1
O6FIra0DTFPCj0c3ImBi0czbPXtJjaciJ8uZlJMWLqoncSEYnrSrLzt4Z4aQCEeI
7b0V4ZqUSWOaLShRraMBjnEJLq8UFSJy9lviRwm0k7bDmBLiHZ5vasmg41zRcaFe
XjQnzE9/V/r6qlaY1P05Y+7YPTEMDHJIbpDmH456jcDk7zUzwbbmb/XIXAX1Hntm
MViEK+pzalkgmS+aV10KzKE3cvUMHfssaNt1E3JCTUXmWa7Nn++dadErEwYVKEF1
CuHGpthO4wdzFYashMdXIrv5txl/OyTBUzd3hPejpQsxuS16TMj/H7sDdSOfv/ka
pPw0o8jxFIw/eVkOSWy9NY1pZT8jY5pGeIKvd73IRtuqUZ8SE7y9AlEQb+80hFk1
fUZyqh/Q+gdC5m0TBidS9e6dwNNcJ3bcUzZ/WIvcyrzlilCtZYnQmKG+hgjExBVM
TaUUM78pBEZXSzbol+nIwKzEPC2CmkKzencqHv7ORjaIQqGJCroM3GfD0BTrrhI/
RKYj+q9UEHkcEurWLfbG46nb0tQqccuhslk9QWcdVZnBrWQXyUkh7M6/JzKponDK
O6k450Fo8WU/R7PJWuZth9mWDTI2X4+ANQHuaP9s13KI0EvRA0xdiaO+VDmJ2t4V
4JLwEEq1xgb91WJeAUC5ldS7aHZo3rojERvK0aSBmmy+rweV81Vushitp2X49Orv
XrtwjiZPFH+ZW74SOXnWnjWpo8ClNNl4bnX5NHdNjj1ChVUWVqxVUYr95sIynuqT
Nr21dwt6lSVLzP5n7/JyV/punq/uBM+WEOnTAxT1NhoF9lgrgj0WOfj9MYQp0C5h
egqR5uYv6Sp7Q/mop/Wqs3gQF9ochEoKatxOrv2xbPtU3RA5pQGwWbWgAioM+ACo
9ImBPCrbl5n91S6gl2vgALbv3yUDrr499DoDHQ4cwzFdlikJgyrIo7VgVCdiRWxm
F7ugq+j0+M00Hivw+mWVaa5qehmtPPlG20cHKCjZKp6dvucIzmJP6CRN0KI0mSWX
4cE4RRLGuzD+BVYkyX1vxP94AQuGt4Tfh2gMcUavUEAkru24Wp407DlS5lChbHW5
3zDEDAX9TwWrg6FiZD/gXrXjBPWPdaF2uyCqZl8pDbjUCHyzLMhc4B0fK101Wuuz
CAIRTBr9UK6QVTVq49C4NnVFwT6TTsAX5MonSbNQKUrZnoG5bo0Ds6+5DbzrUo56
0WgfY4thr/RciNrddDCEj7hYgW5tiDe+T/KbrsgGF8p6tK94HteDm8yoHhZYhRMv
Q/cpKRsZqG6Vn8TyCYnBEWhvezBfLr6pKJJbSoSQrrTio9vtama6YeZVQpM6gbMx
XVBqWHstB50jTvmSjqBxb1XDEcqQxbeJn0xCcXdIVeZB+1PeqLvwOVruBJSH9S39
oGHXtCi9VKSrW7faJ58RIt1o4sQhtjMN7O1O0GRuNLyxy6oYYQVnABbAI1MzhC0u
s/nTS4CsQyAt+SZYZAlSq2/czCOf+nBb+fVemXOcRPj9rbRevpBPhYXPi3fJMg3N
Ojzc3NB0qiTEuLfQdolWjCiPO58qtDFIbj7i0lPHRfl0X7N20jw0A848LXISK2gH
L4AGQ7gdRQv0qKGeU9J09FTWCsCZsnAyAtuM9x7ZJUx/RitrRBevpsCytWRX8oTR
RCQike2HmGpGuKY6vzmvtN7NhjSNMpmxfl3jKWRNe4ecyUZvvLOhYuVlIoFGJTZq
U3522/5vkq0JzUuOYoxAGVuA9YSWAuRolrvCNpQLQ65K3B5NU9MOugjS4Z/Qszl9
I+qseKfQXFKyPbAj1Z7QU4A4tQC2OQ1EHRSS9XULs6AFWekCVIz90cHBCCshsjt9
Zr3ABxjnOo1KjCwefQGEVqr/tyDVzdrA0GxpyzueJ4uxRLrfiU8bFzhcRhXNy59+
jl7hx8tc7rUD0TzwMWi/IKCKpNcv0k2cAvfLEsJRxm5BTBNWW+OLPVd+DuK0m1pv
shiDaRxlYafgmT5dSfhl7QNT5zVIfJdwkfjwPipfIFi/xFcMBuFeK8VWd7hdFRK4
fprBopk8zrGDLEuXma3NNyWJpPk7cT+/CkdMdJNb85/kIFJcko0S3QAxyXq+/e1V
rSdtmCQWC/tM4V3mqODIVYBFdaJwa771bYpAd2guwEcesOsoo8OwE3ZE+hvk8x1t
ivWlc0MPBbsuFqQ41Jmky4zoHtV2NB6RtSElLL7pyzdABmFSPbxFe0WGI1VBEV56
2gVsfZ8luX8Qn0Jn7TDhAWiG6VlOIlaI1u2Je5VmCs6mJ/mH4AiEP9Q5uvsiAW5a
SzajhtWFwAhvON2q+vevTvEXTUBEt4zA0bvOcLMIxi9BPdgvuskZ+wo/Ib7YzErI
kQCdzpiAOumu+D9MkmNk/TpQ2lNoOcSLABYfU5x9WixZkm8TsPSCEXaqMXACYed/
3HK578XTJq5gTbF//7iluY4GtRSqugOV5SPdf6yQPutnzgnm9oDifindxZn2i9d4
bH11NBiYLpdvZ94JfBfPqQpFI7P2o8H5lHpwyCdyQ2XrD/Ff9Mm9DKRuHRoEe3kx
6mob4gE2nUrATpVuOUq92GfeHbFkfzCKRTJOQxowHwCR0cRdOrkqPrE5gOCrIxgc
mkRbWnwI8u4Z7t3mbe+yIZ5nT1k8L/h7/Zapn5rKeVOvujb/VX2BUKT4mhNBoEKv
LFmiqX9XnXjXjm3SHHLXvdobjI3ume8XSeWk5zt5O1QXN5lZcXHDoulBexMSmrgp
eLgUjsK3czUc78On6X22jT8oICvAe3nosiwpxxh8/knLI77001HeV2gGfQhafS3/
RbFFDTqJ7pPTv9WD97s1BnqDKKzzK4JUwsLfqlcy/tOOq+sDs7o7bK+T6efriOrn
BfTr4EIUPqZhh4a2CxbDulTGDaSLgXwe1eXX8mGQgUS5DtBEdFZ+N/5xGNW8Vj13
0hUdDgdPdp8R+rRDarqc6kKlwtY54xyr9A2QBIHsSodvI07YBOXCIZEksSb+bPmG
j7j0VhDsxLpRtaTQPQv71vjk+22BrWMk/38YpvjbAtIPdl68cjxodkWHavLp7chK
+hjNd4AMFCElo501utqWn84qHQX9rpmBR60+NeRGalrWgBkm8KTaBaV/fkFnnYIp
5rUClYLN5VqGEc2pPR8VM+PyhgQM9MptytPlyg8QFHpQeET1yF3zjnxiwzNow66f
qqo5fAytA5gM+wh1Mm2OeDFRdKcKkAjweYrvE5gQrpfcyTmIyIo8X5p3BmPPRT+B
VZotOMkNtQmDct8vCqJMSyjAIjv4egPgpN6HjIfIWDEJXP9GIfVnih/rlAvyw6Up
Bj53WqAD3OUzlLA0Th07KFpWF0oSpdWCmVm9xfkymVWEHQDBpcRp+ZDHz8DV4Wc/
Qpe5r3gmGUKDlCGlIQBWCldwtaP95nHExqCc+C4ApMK95+EO1wBMr3PwjAF1UwRj
qdsBIbSXM0sBTDmdLeb6d1jofYu2sWzQOpYPqbq+2Lp8TKcBJSMky2FK7MnlwIwr
oPVmJ15Rc3rwQF0Vz2Ea9iO8f/olpGx6P08YwidkMgIDA6KcIiu51O2udr1cpKoN
m/hJx4vvmuneyQlS2I8nF8RqCY9mCJI3yfHdVqhO0TCFUcVwAvx6qA2WVp+UTECS
HZxDqFyRVmSvfLNiCZe1VJ/re9vnER1L+AciB0/DgngjxpeliQp2mOGnvCIwwAJt
1Dn/KAJa82gycLILmMOT4FWIH2viKr06xZ7PuLEvPI7DuSvIjuxdlWQgmCXadpWe
t+lKnx5mPUIqtskf0prbXiU5/DTV29Rh1rGR65d0gxh1N6aMFIsPjIAh5IcQ7YSp
z9/bqjOrdyHThUxZj0hYwYe4n4PNKf3MnI5OooKfWF5e2PLRuSYdyuqvcKo1I+XH
Dqkmoa9ecBqYzBQBz4R5hPpQrd8j/pz3Nlwdd4Bhxd2IZI2AmoLCZmdEspzmhzQt
mbthIceKWqmipMUNYcJ6+0cXWGSR9K9aa30sdkxo9CeGM3NY2CIoU9Kksx+bMAeu
LOwB6L1BwIOeZmx6DB8IgmspsT+Fto5rJsYE7du6Z3aRzJy6R/zgtuuwmysVIvJm
UDMxWht+h7mbgxyKg7nNl7oBLMjDEHFV9CmHmnzymj3g/KBChkMmZ2OboixPJ5wj
K3lBWVAZ+3RKbZRiT8poG51fnPWW89jZxSvv+pzOSSWb/ZQ4K3a03HfucP1aOLv/
cepD2onB5Flk4CtpxCNoSqH8a8YXeibvdHeRsBTu+9e6XnxZ8OJ/88S4evSk+3ny
4JZvYUU2hRJ8qqwytcRzPL2b/ARM9KFClu/ntkM5+3kjjv8vHVNjav2TzrP9vVvu
KIFq3G/YFN7FZnWTyHGOM1Ih6H2PedT6AaGuFaghks6UGJ46El0MnfTobPkN2zQq
tS/+jaIhifQkQmRFYEBqIXCdIkNvD9TA60vP5hVyjHJtY3ZQvPpR5b3H0Rmo30cM
O/C/6FeVFBdhZSmk3Rms0ibXpWMnF1clum1JtF7r5WINxC8CI/fBhs/r32BQ5Po4
Wv+KCvf3csHZ9VH3YFgWKWX3Yg1Z3j/og8Ms9WZcqbMpFV1Uoezsyjw/y654/hft
e5beIrmKjo/KFFTvFaZTF9Skcvuy62g5jqZGdfBJqfLENK2QQQHIwAEXmi/KxPxL
VoJhyFBmaPuo+D7j8BvLPC76IYPsvt3oe6F6I8tTbWc99rF/W8ZslXSGuuhuA+EE
cHT2XLnF11Ufu9yhGNngFQB6YKeebSXoWOIHenmAAzxslvfuS0Be+PKRmbmzM3yN
d9Q1hxc8T6Cgb/JSWQB6DwYcgpS+7fLpEy1vBieiMHGScUwvDnCUn4wO4gF0u9h+
mqLhdDBFq8jpUX0YCoGcgLE8+/dUw4siXiQI15n6ARGHUhQWrTj3JEava8PJYOqa
VXPHrIay8tr5bHaYEraoStWZND8H6W7diauOzVH5xVNpWiRqhnuM3+r6L+17VCfD
ZaZJHUb1f0zyQn1UQRANVqrQvinq2UlWpaTLUChn4o5EDG6eAK2OuHI3ptQxuan+
JTis7AljDeowkOEwy4spuF8sb6+7qFSvsSSKddV/Eh6Noj+qqqOUdwnqZD117p32
oWY+ssl6TqynTQGnlAsnpbeBsuVH3RE0cgazTxTGkWNdKnh1gVUSVXVgxwOkv70m
VttG9NMlOLasbEVHPhM8ymqsnwVXZozG0nThfL42ONbiTV8svoayiboaXu0RSoQk
ufKV62s6qXy31mZHOoUjByWMytWNgOeq73z+DyZE/fk6PHnSGJZp0biGRzgTWQyD
wspaEyPSRJ76yQ/0wLjE1X4QH6Juw+2kIvPTHBStJIiiRXmHTV1irsH1vtv9j8Pr
y+ewow0FyMuevgiEGc1ki7rS22dkrgUY8veNJui20uIrK6MwCvHKt0verTXx/RB4
WwRc5jXmywPV88d0mKeTw/zvJKhL3ypCwCR4vKoDhUCIQVkzAt7H2J6t3X+D3Ofd
2wte9vj19+mrpnI7VBojbJxCH1FJAOgykeJrmz8vZ7dATPMuQdH0MmRIoQCMPoG5
gFE63SUBQ+Qhe2aR87IlRzfy3xF8VKhYrAiAezXlUf2XjefmopUKzRkOm7rJBXNe
lEyUFiYkoyuzz5/UJAsYvhOGca3KcQfaE740w38acvhhQwTB+57Qmvd3kvkct4XL
gs2iYNIXapbbBI06IBRLnVtwcUyteE7bTe612agn6WgMBZzLbMhw2/mqJl4NkV7K
zcTs4RiqUO9MYkeUuZNjg6ggOyaCHuHq2VIsfZM3I/LJqZctIFbsKCB8vS3oUHs7
VJrtt3xMbcP6tC822YAZaqOpMBciDLVoVk/jfw3l0ULHSKWCiHr/uAu44wREDCZ6
v7kDmuXSBnc30770psLHI+A8ketjJyjx1PhU6nhrPMwSAy22QaJijU0tA6b76gq5
hIRK65ZacX0r2yIzkrsboWUD4TT3YV2dpCt1PSKxIAPWfV8mcxo3HSZNLsYOZ3Nx
b2KmIvV4f1XnL9W0/ulqGKJoO3D6SFVlrtDUf5ZkR1/TovpYuTJo+AhP8Y/zRLNt
nG6T5MBJKdsmjO8a+Xh4p/0NcR2isP6h4BbrKW8FAG7UMQJEQY1Oc+Y4cs5nBrUD
UECyN7b7J9IIO7rP17FqPtfVa5WMjKGRknIIQHf33MkPqSmzfFZ8TujisDjRpysn
KG3XUPnQPE160hnV3jpk8e5YO+lda+D3mzBWzjyr1BSL1RswWlCMbLHifAeOxdoO
2q8teXbX8v7mhIfGMniVH/1FmJoIN6UaVOHQkKL+Sw+C5zsWoWex5dNQZkqLDG1B
jgy8ikyVHM8s1LXd0mOSeTB+wUgEDEubMwz4K7213knyKFIwTPW4t6Nowaqi6KYc
Th+Qj6dLN84VcS1klwupw8oJ00t1FvNtaM68SULPhemLRXeOaSQ+jN/ZdNgYOthy
M4YqMDXD8pyby6b0d0EWU8p05N2a3jKR0FjiHaip3YJ/4rgx9RaW0FLOMVbWW6W1
NSONKU2DDZOpvdLPHVogL0W37AiM25r1Py7zKzS1Svdb7hYfxM8W033FRVGZEvzy
Z/N2+YT1G6qh+YZ+XHu2LaBOMu9++xlOx+82LiXRqiK5/AvTKVc5u7uSOiWZkYcO
zQbycCUOpG09VCk/jsUFQBzekASUdsbhLERqINPhptPLyZ9ruO/ZJiZBj4tsCGST
eI4LFOjvw/6wCw3J6iYxGzYq9fDRL0eQl6ticcfaFTN8P/4CirQrlxdUKbe8RdY+
pyF4m2cTdMgr+7EYedUYOeAUqQuaBYO3S00oTyoX4uKqFeTVRx5MNE+uQ6RpT4zN
AH1UWNjyyn8AVmm3pYdMI3yzsuxPcE9XRtywORHpyR4scPGcOnZkhF/z3QZIkwgy
3EGoQuuh/R5rMEy9ic7m/0cXMVpV/BZFDn0df1ZqKWoVIFm6bb284UzkilF9ZUsP
H66rSkVHj3/Hv6UlAoC8iQj2L5j5K77ER7BXs+CH1tjSlAMvQTL2s2CPhZavOYS1
OE5T8/xOQ1iLQb1vMuff8INcDgPpCNjkB0fLSU8ibLDTORAntdtbMWVthlSggvzT
BTzS6NJCPEBDCCZKkeczHvDFvWh3/GMrmxM+n1iz6pw42lwFoI1uxyrEyMU2l/Kb
KxRvkfpy6mQ4eyi6f00IrGnFDACr89mIp0ocIV342j0dzzVOAhT6nMoubKpbEIbI
jTkJAlFUOb9MEe++g9AEtHRAOvym2JfDzomzmvoxyeff50EHM9ZFe8Ags0fim5QB
gxO/g73Zk0Thf6MdLufyo7Zt9oyAvr0+rOxKKehR3OMDgZLGoldnTAIHttI38+hb
MTq03G6suO5bfnto2JEtMDxhsAGFHSKd8uSdirmUTZAoGnWwZSpVWyMScK+rEJe/
YcU/8mjWkC4+druOzpLHXzIOHseytWJJ6wTx8uUx+gPV7KmoK2WHrciXXJFtLxbr
2z4kEaiY5kk9JgQEfUPAv1botZD8z1d4irTUad28NFmjsf3WLJUgEtVuTVgteAYv
lneaZhpv7WzNS6M7Y02lOja3UY9enamV5lDwI46TMNgcRLTybh4wdBYChSz9E0Ki
rgUOr7SGPy42/Ys4NFheaHSMj75QuswDXIMj4JRMpTeY/pFCfjt+RXdfwz6KNfTg
7UGDL0xzn/1LFFIhukneLCw1qJ2rQkA3T8bK1EAq3jeE+cvultWmA8PH7hUNOY6l
DJnOo9zSfVgRR8i7LD3NlmiKOgYK1voduyAqjpEM1qruxEiUTVkHCYmSFjLeAvd9
ZnzrxnsvG2c3fI3beR1lkD6kPWAhSBTleTbTicIOpalQ4DfHW0+nyKvbhOkQrz5b
8nLYrX1xYPDjbiNRlyeTt/A9CnBk+hGJsIq9jyM7LDVORbiF2zdDRqCXkOV9/p9i
cdorb26cZhOdPKk8Atr6VH3WP5+rU+Q6uDPGGOhSpEkdWAKcb7QxpwxbXo2JwCWQ
swiQlEvN9lpysczteKXYCV07EtTAjQ4TcO2YSyPrEdAsv6HtHTjdr7Z6nS7DymoU
tLgbW1IYFG6MLVhQaZqcOylnE5tRHQD7TqIx28Ea2poMfmm2M7HEhf9Bd7WwT6Pb
pMgXRgHjBYpyYqQn3iNDIJAg79WOJo+B/+2Ee8UEk0/k3VsqBg1+Fj7W92We9aWd
5nO978X29SifDtPYynX79FwF3iRHp1Xd0+7VKaLaJxKuARfysZcR/T701KDDAFL8
XTRTmcRUYjTHpuBho39r6XMheWlYff0voImadO0859QZsi+iCCbICpgLtklUXmKS
pYTg04uTUM09KUB4RBT7vhSSsTTzlRrWkU6JnejPH53DyTLYpbUfMtmQNCC9g3ye
d/lJVRNQKmTNIOaLQ/ccyy8THqAMj/kqKAsBfHGhLgSinEvIkxio9a/Abjc2QCZi
X6AKIyFCQ94aRWkTLkBG+zZcTrs7HPhotwHwFmq1b3/PvRUxvmXcximvVzfIJE6Y
8NfCzgaXdN70nHSw/a1u0pBytxjfUkBzjS9O+eHxY5wP4nnAz28aXUEj+Rzxb7xV
471eKg92MYlVkDcE0IDhRE+Ixqm5aiUbwKX5SFhg7ippPCpDO7ysCxsXSLbX+XTF
zZUsw5/k5GyV7dJaB3kBavwmlBNPQuwxl2uqeEQoCrQ5jU6pbPOHpVQTC4/saKAF
TxxBDmKfqUKMN4+Qmo186aLOcLvogvupJTSMBssII2D3ZOT7vLAdHOFNCsq+v8io
gszPW1r4VZxTgcnfIV5aE0Ktu9h//3yv+Kyd8N/cVYyEccfF62lzuc0jtXzZOJyM
p/0rkN3ns2vmo6PYFaTTNlElWymaVaOlUIKjb1loPdNuU9dwTWAiBanGddDVZNEy
WD1ejyhCchftV+BfEt5fWM58UTW1ZPUoxNWYuBBARVxgb8tCWOUDPqeZezQdZIHe
eZZfphbEFj3PVC43sXIRtGvnYmXKlHnDrSVlTbm/nH7hdm24fyfo6y1Iz69+UHV3
ZZIR+6Ly8TNCe242E4T5Ayhlgb4TYvdf8F2KiUEl90RZT4/+B3pjj5DehyqFfLrL
vP0eOtaUHRzkZtKP7kJnFTxaFBcW5sPpZLIEpCmDl6ORGaIdH+uYQkp9E3vUCVZw
sP9WX1jRj83egVXFtJmV2799voG7S9SwzZx0zA8sNkmtHeK8NDHkI/NrUgYI/P/l
affqz37jQyiTjxrR0ODLkXmIcI9ec+dUNJqXHgTfR3d9HxL5OUKhqi9kFSTECrar
aIlwRelIsV8xwdTbAtH+YbDMpRUK9cV1okOloJ5UJCJ7W8mEHSMQ9TglKYeTV8VM
yizGBHI0kG5ULE5dhQ6wYf4VeeY1vXBsQBOw3w3OkocLVUSdgWH6pGhZEPTAo3gp
04qqxONLS+fLvalbBpU1x/PLgfwfQOIoZzvc9edymRImE0+9XSRnxWUZ7+iC8LEg
xbBVRX6/usQiQtHlnVgV+AN8uHnY12MdlN8W5Sk85QI8t6aoWD9KDVubWCbKqfVm
e7A8re0mqK+sXqPAvH+cn3gSwib2lCcvuGo2Z8cX61ca6NBGNJZKQLGA0lIMv5th
/Bfsgwy66uK3g5ZiJ2qsrA7rHPn5MCTNPxtjTC+JHzcw7flAqpJYynnsfGug6GzW
BxiGMxg5DN2yGTmnCxru5T7GzH/svF9hhqr4DvCNnOXEiTVZvWHoHtNyJWrf+8aJ
ChVfG9j0bkuwiwIBdEjsk6sIaJKnndIZBtNAGpHsKtG9HhjKLKmm9u8ryTg1a4yz
x/T2J6MML2tJqFnFZ4+Kzkac2RYMmiS8L9D4yYprXM/0RXCK3sgoTRlRa6v4tPbU
KI1d6qPh5z3vhU5kHB+G08bU2fOLbW5LXtIbN2EpAeyjhYypRyZOhLDFD0XNvsW2
F5DMukr5F2qIdopqvf5SE/nuBi0HzToXeDDXm/UwqxK+b38ccdaLJWJRjQGh7J3l
Kqlelw/j+GxhqCvxXIbW3KuwHrqj0hScrVsBI6wXCqHwYVYPlOizCb/SCPqgyTTT
3/hYgF3w4GYI6sJ54LKh6hgxHEGhd7AjKgG14QlNDVDh0wy70zdWttOeKd/j9YcN
r1N7Pf6tsxDYJNNMxxbxjPh53T7nr+UIoLb3eQMmJTu+SxE5u2Mnj5L3+Nn1umRY
g+5psz9f70mXzpPgzHgM6dbcTKmyLrENwql1eIa8/BD1MHWS1xBgxlCbNiDidFSc
iaW+o6Q8EYhwNhyNunRWdQFu+ebsFzP2JMejqmj6vLBG0rNOuTspoE1M4lr1bA9j
7OMYb9YWWqlNSdeitMe+H98k3cv8yV3ApGXb4CUjYxtEOw8uarjQp4LhXmuzlsok
7q4nAWF0aH3ZYz7oPXDS/N0JaHMZK2q/9Hpp0lrix8p7/dmUMtin93oBZVdEJZ5+
v+oEgspx3IRCY9CN6a+MEB/EI3HQei8ymmT2qdPXVAb1eMcEERzMP0c00euseBbR
CNAhIWOSz/BR+paP82czXgEhuaZOum/gKIGQ0oi6pZ7jTg0rURX94Y4kIqVPw6TK
GlgeGWhrq0E9x/ldxvImwC2x7XUQmfT7E8zW1Us74nYHHYmPLG9ofjgHl21nk97C
ZwhsBvAxL66a4+UcCCmAEktIjG6W89CoXOL0kal/jxnym2kyBIv9KKMmH7WulzgO
L5Dft0RYyHrmtb8HAAmsUWMy/B1PcmH3A5VqBeMy23hG3mVlvl+8Z5eBI/GI6kjB
sqOb8tmaHUkXmq88TiDdNBv8+q/qOIx+kBXpc855w6sbXKGprLnTttaV+Slz/RYs
StdwUgI04EIAhNo/Sw1jKrslZR7lrY5BnIS9xcx45fplwgx7+5TBb9J4MGYJEN3/
0UoEYIjcHx6thMCaXcKg2NflNGN7mvjyPLjKCxZwIIEbkzXeyFIeIMemiGKaKhJh
mMkXYcvDnzF3K0bAXX3eHnkM3wS8bigO1dk2f4q1ZpaGMGs0QtLLG7/7ie0Qs0WE
ul50oYQPvlm0+ueu71Ljr+2C5/H2LzcrvNc2G//nFdzgkP22qUw53cF5++0KJmWo
8PC7UNBvvwzp6h6/58q6N/1yBwWzYNB+rSbGBSb7lx3E4sQVje74KSzS7ftrxSI4
JMAI8mJyzM1+/T9Y3V9+U2NjMZou0wTIMXC4cBQS1JNOjh9dQ16y3hYkz+hP+9cD
nhn4P+qqzbuskUJPMuCTzIfemI75y8FKZuyjy7jeuOJZyZs79XtnxmnL9OMIWP93
4+VwEtgZzhK0Arp3RKGWUVMDrUzBUe09lEk2BawjG9MQx6uBT69baG8L7cbe2GaE
Eb7DpImJQlIIqzyZj1T7KcGtLnq96Wrf6MOo4zGwfd0ZlWouMmm2kga1+blv6dj/
aP351X2DdkIQ3EnZKGLWD2ORWBP+3drbisLk+DSHe6skS7n9mw+Cm62TnMWshi6F
q3223lV1iTS4XQhsLbbr52rC+1CgVElCknV74fEYc74f3rD6Hgv+KGEeaeEpKhVv
Pewp4nZ4nAZ/tYV/qIiaAljehVQjtTkogMTwrjifejfcB3O/+wCTyp7bIK3MoDQW
ZYtfjvkZaWL5F5zDjtAw95mcwa0rJ1gcia0mtYS/55UaBpEYG45weGwfYxTxh0df
tOC1WI3oR5fdtl1sHTE6pGcyyCa3Hfo+zpxA+Ao6N3Ridw5nZ+KvG9ls2hwqDpkp
ZX0KbeB/geJ6JOyU/bKfsm+17usMAvWmHMGb4EBvZf+s38Jn+nF3/Z7frHvmOH66
h3WkvM2tbrPEiYfjxz0zZR/bP5i5XNegkn0gvH5UhTcFXWCoqjQhtGLjMKxbWTFr
8YtklKBtGdcN3t9+qY43As18vbNMJZUplyDCFR2MDdfrRyYwyz23OwCWCwIgrvgJ
2EupTS+NR+onP7sEbhkL9BYisxaNDy3dH+Vith0OobOdJfQtfqYYt5pJnuG9FMHB
H2owd1awdFrCo5CoYzoEdwZsy1pYSQDfMLEcNAG91U7/72We4MRp+UTc0L9xWSZJ
r/kcIplZYNDOu8qysILd7v8VooFnWRw/r4Q0IkPVFLEZGk4aM3hi1tl0HgWeON45
B1AmppNVUMUFsIinRU8wFY902snWZ4HSPBlp8TfC4K1U0J+L74Mrnd5xzml7BFWH
Kt3A1CgLPtjzEeBT54wvPcOUXijz/j3ZcOdLV/6HK/++prLtPEG0x9rC4iufyP3y
dWLT3nuQcbLCgY9ErU30eFfi2lXOISWJap//lum11Md0YQufAiSxEeQJY3juz9Gt
5kdWwMlsQt/WHyIKI4X+7krx6bNLitw8OI5djiAPiULeZnKBshw7Uu0HJ/bkIAeW
6Pp4jJcXTaAXJ0OyX4zk98xOTi6BE+i/XX+dRCEYLGRn3Bcu9huS0J07LyNTGc+d
W0GUPPtIHFoNVDNTWO+XJu59qLmcTYMUx4aHgV9pignki9EJq0CwJWXBhYAPXMzi
Q4XuQy2l0WYa5HPClH+fYj1SlqayfWMpHkS60T8/sRRkYT6SoCX5mP5Tx8XnSVrp
gfyxLb/3jS8ukrpvie1qJRnfbMYdtTHkIFORVNcryOwcDEekG42C7Av/7iFDyhcx
kkdYHq48eFpYKfLwsqh87B41orKubNqBB6gLLT9RAbriHQ7Gx+EBV8bEP/QsU6rm
vIqKWxi63nbVggFiN5XSQ/lSiN7I1Hw3O5PbXq9V9oIdDXT+Egn/bO5gtEtVlxYu
A2X06Lwej728ucb89QzksiO4DIsNvIbcp++2LMLNkggHrX9XHb6ab7YGSfeYfjOT
HF3yDmB4ybioz8CJ+W+7OjAqim4cFoQmWPM0zoWnAIahi+sg0ShdDDZhE5+ecx42
fKB5bjD12t7t7L2oSdwEOVnSDkFxeEyaSB8QK/xZnE+0G/a7X28Vt48v/UfsOI3j
EPOSvA/q7uRLiMzqZ7cdYamIOU6tCnsdpx0ZMnGzIEycCrMhlbtBJ1u39yvTlVhN
cAGVbvBKKUT9vU8SSBZOFPUtUPUd8yMuqc82TsKulziyYW1OVK5zH4yo5XIPZREJ
jDOWEmWIjOrBeOHmNxnxUI+1uhjXBpyJhLMLFZNPefOxh8dXUr1SL+OrRIQ+BUip
fb1B0iGHKxlqhGqHOLJDnZ74xogfOKKGQpczGfWdOQ/020XjUJEtaaSJA50rqxbt
9e8JziDjgmusLuVfsVvKW/uNXD5FdG0uvDnbpcfgC51VkEKP9Hyv86mwekHfINMK
OKDFzIbJq9RMEKVwVLlkfre07EcsuFQGcrSEgLwFXmSFmYDek3M9C9VGsqrgka75
mqwe0FwQxap5yRTpoEOKnBc4eKxa2h5Vh5UDK/xkzZ++GqOmnq9jRV0LB7Kn19IV
s2WvvKWLxyrtYMhY0HVQFX+UJpX62AD2RXEojjq+Fi1QZQ/+O+5qfy06HekPNTJA
URZOj3fMU8W8BNllZWp+tSQgQW+GHcKigjempgNSKShenwSy/MxnzABzwHwxMh2W
eukFkGkt/uETHAmnZNtX/V6aAgIJ+7CKmxESRgG/G9sjGhAn5pn8Wqj6DvYG0Crb
//JteYwYwunKfrj+zcDpbMUsZN+Y71qmRYURgkuYIDhYRDHjjY24bhbOUMOKwvi2
6Oz1YLizaIG8pUZaifNU6GjNxadGKpSHuilwegn4O7Alp0R5DRN1KVOLWWiTjpRB
qthX2zBz8oEYvkDcfpDi/7NEYA2BSuAsWl5yyfO3HqDJnYjBe4VouqEROfowtZuo
n+1fegVrsmEESjoREyWkPF6UQn5vK32UMk9S3xhnG47Xrszw3HGMoskeD2e721GM
Zc5gbH0mxsoHPd74H59Y/3J2ak/xyYhtdGl2yooSBnzkkYKayjoPTogTXyod+hWn
kAlLWeOcIGGAvEHOiBohoGatZoWr4iNDO/pep7LBfw/J33+90O+J8FWPAzR4qR0K
6YFcvrBtyFVTu5gnHXSP2MZ9IfeMBn1EUIizWFpp+tYubED5D6dHjwWMpOwXX+Df
I8v1sdj087taH05P8qGLx5DbuikEU6c1dD4L/HenzjkYtinu67YhqFQCsWv5Wp6u
rrcHsQcxYlgA6nr7vWXkOuMmaD3S3/wx9Pc8HhRW1yaRwC4E4ZcE+MVB0vM9100G
QXW05jAk9MrTvn0tYNiddkqXZkVcY2gBcsdL/Nj8Fopb9/YmHEXmXVh2urJT1AdB
SYPCDYFfjK0j6xQ79SiLYDqsDHc+O+EK1tR4gUmfBZTb5TA2tfVVTk+tzhXprjcF
+WHS7uuQqzag9K76NKxPVbIJkGwou2xcYoYYWvbMhYpHIS7TG7FLORposHqFFxAZ
60OZUgmjoZHSmoQ3zF/BmTuGKxe6iBDohf7YSoNDPRQgvXEM2EyXdYP+nXEZQCMs
qjwwGBcGO50XJV73m5fo7Gq5/p321rTPPa/Tu43GHHKJTSPt8Zxzf32vdobszF1A
ZYA3JleZzR3rDY76twoTojLR5A3EZibop3kN+a5iiydDUyZYEpF5C6LH2ZbB8UI1
vs525OZfFcplpeiw2jmSdJOT5Zq5FFc4uXMA0coqU6ggrfsWKVGE299gpEF5rnnX
DEdx8wmgp4bbTwS6GpOJAVCxFlpQ7t10GLFJnnqxz+vynptuxoUM94Q7asirbGm+
rNKUNPaWXGcFR4kCmor8875KTpAO0Ex7gpIpxYmRGfyATIWN6TTThsvn5ukE5Qbt
DbZij22E51IOQ0B8PQwKiVmdpY9m39Lo6ZLbeBvU4YsHtzfAL/QdMvGbPhRYdwBG
VlpOIQuPW6NtPRufNnHu4STiBn8k39XaB36sjmGoJx3L01mYqm9pO4/J6fiatkFF
pdzj858pa40N/CBUBa3ugesLKVJbWPt2XFDwI++c32jd4zIS3Tb5kC3K+8/7rvGN
4GeFZanG/1DZ/sVlrLMawCkA6eLo/Na1iQ1F30d2YudtD6fKCUEPNaIUuXpKh22U
21Rc0BT8QjyF7HGcvD3GlufYwRHLz4IgKNhDpvJccccXCSf2ISuuj8IKLO28cEmK
jrg4YTlavPzP/EVAyg92PY1cs+yb1RuFvZSfeo4WzT2kLAMdcq9/USMkOuxBpW11
qSp4vJ316TBGMOJvH+fsI7cC9UMjYXfyLz4U4OY6wOBEwLDM1bpCScJgNNHzJyCW
gJHoadhXVQJEXC3brNhkWuwquogi7ZvOWG+xakbsVuMZWYlMjlZ1yBy3nbCq5H5G
zBWWDmWJX1E7W/bIj9XYpmnaqk3GPf7yG6Lk2CGtcif5ieaDfcwHpK3LXiqkvdwk
K+RXcjBxxb1LrdpDYlfLTG1/NqLNAxJxdUVm60JUOdkz5pqmHS+wdIkkNqH8Z9i8
5XgXS5KPZO1+/s/J6fiirUwb+rsjM7TmIWkFU/a9bcFlOY7GKEyLgOQkMa7lJ6Ik
4eHrL1jiFnhKkW4VwuUSctM/6V8inaQWk0grelCEp05sVKrLkDknpsNv5J0sD4m4
G6meWH2q3/BAo7gx8KxtIX8Cfqvz81vWCPqf7k+9phMATS1zCMFE9jQgSx12sBEp
667jV5H+yEYis93f8T1LkybBm9feBRxN+uVsGdKR8zTUaVzim+wX9iyxJ6YxCQnG
yP0kRnmQKpUkNlTp1SJZwFAP8Zap/3O/kdxTJgr+v+LtBk893QOYGPUGUUk9bV/2
qmOTrNX13R6hFKKYcim44pvhH8tFiPjQeccNCOrNeLYvuiEXlsn9ZobL0Ke8lsAM
ntMT46D6hBYdOBMZ9rFQSry38rB66pFrJUVpMt0KoMQ9aMtVc1+VSoY39WZi9Syz
J6nPax4WTBKBolsWQuEFYO3aEuxpWsErgRBrJm9wMU0H5lrs8gNNs/qXeIKA8fqb
wDE564sbAcShgSVPnpmgWcR6fNwvnYtP1QrQvbmi0SeTQxleC3WDvStMEFrEli6q
7WOrQjWebbQ3xwFFF0qwW4o6cfzJZejJO5f4lzksg/v9uVl33MjPvIj66SUgf885
MUM4B0Y7iHN+Fz82hHDuE2MfVMJHkikHFQgkk8TFt/X+X18xxST3dj6EGZXF78LQ
wFovHAf9sfdwSH/2QR6rltAZL47NHNLubavvfvf/5mxglTRVyKor8IlNjvvfyBlZ
MsFT4+np7W2WbVz8MTK/mXT3iBfHfeZwdcfFSvf5Jyyd7+IXfzPnl5dCKQBkNSKU
AVOBvFqvuzDlKOTq0UaWTSFOKDcuevNpcdj+GdQpBvEr6MkWyA00GyaT6sI8kjQK
8ftKLB9MVK8SJO7g3Rv3RKoj8FSOgGOeRngoLR3u4DKsS/IAtnHkoFMz7/Mcg8r4
YtzmXphRWcUQSokH6NeTKbNKJDA2X2RxHoB2TMep9RCaDmhRzL2ORJPlD08k+K3k
PPI/T+gdIiwrbSoPPd2hk0f/FqRwqF0cmnIbs3G3na/MmmdTIhTGmczM9A34gVtS
o1Azkn50ZPdr5pSvhCwO5XjiOQBgdahqfRv9gJhxNP1ULdADMR77Z09nvGbxo26y
nZJmhpxmG7wfa2UiUumgGjkde4a/qsEpJ0WTeGyG8eERT6/xJgKddszRDvdtAJwt
0UXHyxqQSe5f6L6SdBHwXbjTLh21hW5WSPJqq8OHAbxSHQcqbT2pOBkgiBcdoQ4r
gaosePcL6zcsH0WY1vvrYxvyGSQRfXYtfHA2xvFILK8NhALFBBG8vpSAsHid2K9V
QWSiGLElUlWAg7f2ZXFxpEydp5L6xzOaaid7WlfvgHIjPNu9pj0hTSHJiQDcUMf/
GTOu64GeRo2JWM+mGAN9JO/hoE1J/cr9I4xLX0mWfNG7eQikSlHFhBm6pXwde3Ty
aMhgdxu+Z6+gZbkbVztmLEw8o7qmrUvfjV6pdBU7P2WXptxhYuetTiSRh6irugxn
/lKda2JZBR8XRWq42W14y/AEF1j5cmyWECGWroQRV4QpX4HlTTWYza3EUCG3DIYi
HnNs+qkNbyZUJdamTFKHXhNM85PY6kKwx18mafO/HYSsAzOi47yVVWdWralKsDr9
8OVZ2FRlY7q+XYex4maY2rMZ/bqprW65sOffEMK08xkrFzFh6j5t37n/2By9Qcqz
MagtZJxz6GACJDAs/dKrDWTLuFj2RZ5NB1SWO3Xyv1Tt8SoumfZO2YShDz0RuOSd
9G9ti7Rsgmi1pXv1ClexZGDRTPgnN/ultGE+7Upq8RjqnpBpX8fhkN6CwpXwYeEN
eZ40ump2aqnHtVvbf7iRTivn6Ri1CPlPPVKSxBP2nzM6F7LmqLcO6/c8LiDqV2jr
e7HtVPkC8anyElCYsZLJLlmZodYWYeEfq91zsKACiD+0+KFP0N2mX4U5ono7dR7p
IaCo2UQRHUMu6zd7pTYHr/xPslpUkZgcebWGVdYzQumMMny8QznwqeePedQuNeHP
UUMtl9xaxEP/s+Z+PtochGwTP95b7+SsVUqP4d1vISm7FcDWaNKjKX0aEg7RJHfr
jieCUD7vTeouqVvmBp6z7LucmCcAbOeuTFdmkXy6x/qkR0Y82+rFUufGMxoZ01Sj
qwy14H9sgvIaYf5EZePq/BUBozQjUFPajdgcIqVw/lCk5+NKoebC6xDeuCuDO9ca
+STdqbyae5S5ge0SV1S9TxFYaK0vfvLjAe0O1nnNyQTEDZAZTf82+tkewjHUb80G
zW2ZI0//lRWBKrLlcc585s6c64pUzHEyei1pNGjj9IBKTsjXURRP3UXUivsA/9VL
lpPYFusiBfaN2HFc8xGuAqa6TUlY/0RWWfsh4iwKiST9pGW8N981SZjDxPNEcJ1W
60NEO/7+LwBrPkE/yLNE2Hg/bJ1vBj1gwoIXi0Z1co1HI4U2CoFYINZOdftcx5gk
jWVrYfDL9eWoANBI5I/gpHkvo2UaVqK5oA6l1GKh+uzR/kOTqZKdy4y+JEOPe3DP
vfggK5uNMEnRmxciwDiWesqT6rSZZyxLIGH2SnC2RUTldj+CtJpIqH2wXKnp+St2
SD3K9kYlRzYH1bQLjICjYDuQ/97aNpwyJ7awwCRBBfieWG6l9McS+HY3TNGVzqrK
oZDXT0dFPgBiWXpWA+rgW/tkAivIeGE7DgPHtI0BJK7AfZNpha3+88lmnY0Yx8tA
C8gAZmmqIdgjcFtp1WJ8VB6jkaC9sgHFseh7mNk2levyo52J+OA08MnHp9hwWw76
DK6yfAji6+RAzI/MXrRGP/K8z5qy2QZAjmQ/oN9BEyOEnNFyY1fgsduR0wKMS/xt
6LQAuwwGJrR9RUwOXRquPtz4D4Kvrw8+FIt1CGS8Viv5v6JKfldY4UOt85u5C+/Z
Jo86uzau1nIEDw3a7wycUABqsb3Y1nxJqR947kBfeXDSwqC32k7pyid7UhgYVhNr
NX72TxC8bCsVas1iA7FnZOzsmuoU9eoriqwoU9mGdhqJPUBWdjP9O9uJHiPucCxi
/dB0c1Ql5f/2+4CyZ2huA4lBdL3/fo8qA7KMBdycNB4JVF5qGxnMwT9xyKjuTMt6
3c+ZbNLGfla3MHqvLFdO7b6kfppfin/4Gsqhr78OOtyVejJ0q2XiK7nk6A30SjFg
duzbjpf+WjsDDkAe2r7Lz18hwMw9yZNsQejH+5b+05U1ABN667UJgexd2YZuo32R
FXRiy90LhGfP6mLPGFb4XiEhzqqiAu6H+mIkPVrrDhdi2+FHn+fyNT1HPF0jHcb9
bqOtpCoI1nZKPtdhC2JCAe+PWztZW9z3pSjttf3BQu1p7yJhHEZ6gia8Ng7M3Cb/
TCHnxFiEMlcikC72x4laMCa6fjddI3cNbUK32k0iLMgP2TPAJlbvtL4PU/auS4eN
6GEKx9H0uYS5AsnSLHVWmHWa6dlClvKT9pLNinEwZi5NrU8K9DLouQWmG3lykBTO
Mon9gVIv0L7FEDE81RnDH92I18QrcP1TmNMKhLZu69bDPZQ3Fs6SLs1kS4me6Yp2
FtwRr70SDLaWlwgZPX0hiXbG4aykxeRkOZ7iCBNyGMs=
//pragma protect end_data_block
//pragma protect digest_block
NbdRLTRLtLek+vF4oCRjhihjlKI=
//pragma protect end_digest_block
//pragma protect end_protected
